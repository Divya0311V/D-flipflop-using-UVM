interface dff_interf(input logic clk) ; 
  //signals
  logic rst;
  logic din;
  logic dout;
endinterface
